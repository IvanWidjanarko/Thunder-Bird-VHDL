LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Thunder_Bird IS
	PORT
	(
		CLOCK, LEFT_SIGN, RIGHT_SIGN, HAZZARD_SIGN			:	IN		BIT;
		LEFT_C, LEFT_B, LEFT_A, RIGHT_A, RIGHT_B, RIGHT_C	:	OUT	BIT
	);
END Thunder_Bird;

ARCHITECTURE Tail_Light_Controller of Thunder_Bird IS

TYPE		STATE_TYPE IS (IDLE,LEFT_1,LEFT_2,LEFT_3,RIGHT_1,RIGHT_2,RIGHT_3,L_R_3);
SIGNAL	CURRENT_STATE,NEXT_STATE : STATE_TYPE;

BEGIN

-- Flip-Flop
	FF  : PROCESS
	BEGIN
		WAIT	UNTIL	CLOCK='1'	AND	CLOCK'event;
		CURRENT_STATE	<=	NEXT_STATE;
	END PROCESS FF;

-- Next State
	NS : PROCESS	(CURRENT_STATE,LEFT_SIGN,RIGHT_SIGN,HAZZARD_SIGN)
	BEGIN
		CASE CURRENT_STATE IS
			WHEN	IDLE		=>	IF		(HAZZARD_SIGN='1' OR (LEFT_SIGN='1' AND RIGHT_SIGN='1'))	THEN	NEXT_STATE <= L_R_3;
									ELSIF	(HAZZARD_SIGN='0' AND LEFT_SIGN='0' AND RIGHT_SIGN='1')	THEN	NEXT_STATE <= RIGHT_1;
									ELSIF	(HAZZARD_SIGN='0' AND LEFT_SIGN='1' AND RIGHT_SIGN='0')	THEN	NEXT_STATE <= LEFT_1;
									ELSE	NEXT_STATE <= IDLE;
									END IF;
			WHEN	LEFT_1	=>	IF		(HAZZARD_SIGN='1')	THEN	NEXT_STATE	<=	L_R_3;
									ELSE	NEXT_STATE <= LEFT_2;
									END IF;
			WHEN	LEFT_2	=>	IF		(HAZZARD_SIGN='1')	THEN	NEXT_STATE	<=	L_R_3;
									ELSE	NEXT_STATE <= LEFT_3;
									END IF;
			WHEN	LEFT_3	=>	NEXT_STATE	<=	IDLE;
			
			WHEN	RIGHT_1	=>	IF		(HAZZARD_SIGN='1')	THEN	NEXT_STATE	<=	L_R_3;
									ELSE	NEXT_STATE <= RIGHT_2;
									END IF;
			WHEN	RIGHT_2	=>	IF		(HAZZARD_SIGN='1')	THEN	NEXT_STATE	<=	L_R_3;
									ELSE	NEXT_STATE <= RIGHT_3;
									END IF;
			WHEN	RIGHT_3	=>	NEXT_STATE	<=	IDLE;
			
			WHEN	L_R_3		=>	NEXT_STATE	<=	IDLE;
		END CASE;
	END PROCESS NS;

-- Output
	O : PROCESS (CURRENT_STATE)
	BEGIN
		CASE CURRENT_STATE IS
			WHEN	IDLE		=>	LEFT_C<='0';	LEFT_B<='0';	LEFT_A<='0';	RIGHT_A<='0';	RIGHT_B<='0';	RIGHT_C<='0';
			WHEN	LEFT_1	=>	LEFT_C<='0';	LEFT_B<='0';	LEFT_A<='1';	RIGHT_A<='0';	RIGHT_B<='0';	RIGHT_C<='0';
			WHEN	LEFT_2	=>	LEFT_C<='0';	LEFT_B<='1';	LEFT_A<='1';	RIGHT_A<='0';	RIGHT_B<='0';	RIGHT_C<='0';
			WHEN	LEFT_3	=>	LEFT_C<='1';	LEFT_B<='1';	LEFT_A<='1';	RIGHT_A<='0';	RIGHT_B<='0';	RIGHT_C<='0';
			WHEN	RIGHT_1	=>	LEFT_C<='0';	LEFT_B<='0';	LEFT_A<='0';	RIGHT_A<='1';	RIGHT_B<='0';	RIGHT_C<='0';
			WHEN	RIGHT_2	=>	LEFT_C<='0';	LEFT_B<='0';	LEFT_A<='0';	RIGHT_A<='1';	RIGHT_B<='1';	RIGHT_C<='0';
			WHEN	RIGHT_3	=>	LEFT_C<='0';	LEFT_B<='0';	LEFT_A<='0';	RIGHT_A<='1';	RIGHT_B<='1';	RIGHT_C<='1';
			WHEN	L_R_3		=>	LEFT_C<='1';	LEFT_B<='1';	LEFT_A<='1';	RIGHT_A<='1';	RIGHT_B<='1';	RIGHT_C<='1';
		END CASE;
	END PROCESS O;
	
END Tail_Light_Controller;